--------------------------------------------------------------------------------
--
-- File: DualAuroraUsrpRio.vhd
-- Author: National Instruments
-- Original Project: UsrpRio Aurora CLIP
-- Date: 19 July 2016
--
--------------------------------------------------------------------------------
-- (c) 2016 Copyright National Instruments Corporation
-- All Rights Reserved
-- National Instruments Internal Information
--------------------------------------------------------------------------------
--
-- Purpose:
--
-- This is an example Component-Level IP (CLIP) that instantiates two
-- Aurora x1 lane cores that run at 10.3125Gbps on the USRP RIO. The following
-- code combines suggestions from the Xilinx Product User Guide (PG074) v11.1,
-- and implementations from an Aurora Core 64B/66B example
-- generated by Vivado 2015.4.
--
-- The clocks produced by this CLIP are:
-- Port0UserClk: 161.1328125MHz
-- Port1UserClk: 161.1328125MHz
--
-- The clocks that must be driven to this CLIP from LabVIEW are:
-- DerivedClk50 : 50MHz
-- Lite_AXI_AClk: 50MHz
--
--------------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library work;

--synthesis translate_off
library unisim;
  use unisim.vcomponents.all;
--synthesis translate_on

entity DualAuroraUsrpRio is
  port(

    ----------------------------------------------------------------------------
    -- Socketed CLIP Signals
    ----------------------------------------------------------------------------
    -- This collection of signals is REQUIRED to enable the FPGA's IO ports to
    -- properly interface with the 10 Gigabit SFP+ channels
    ----------------------------------------------------------------------------

    -- Multi-Gigabit Transceiver(MGT) reference clock differential input signals
    MGT_RefClk156p25MHz_p         : in    std_logic;
    MGT_RefClk156p25MHz_n         : in    std_logic;

    -- 1 Gb MGT Reference Clock
    MGT_RefClk125MHz_p            : in    std_logic;
    MGT_RefClk125MHz_n            : in    std_logic;

    -- CPRI 'Clean' Clock from the LMK
    MGT_CpriRefClk_p              : in    std_logic;
    MGT_CpriRefClk_n              : in    std_logic;

    -- Recovered CPRI Clock to the LMK
    CPRI_RecoveredClkOut_p        : out   std_logic;
    CPRI_RecoveredClkOut_n        : out   std_logic;

    -- MGT TX/RX differential signals
    Port0_TX_p                    : out   std_logic;
    Port0_TX_n                    : out   std_logic;
    Port0_RX_p                    : in    std_logic;
    Port0_RX_n                    : in    std_logic;

    Port1_TX_p                    : out   std_logic;
    Port1_TX_n                    : out   std_logic;
    Port1_RX_p                    : in    std_logic;
    Port1_RX_n                    : in    std_logic;

    -- I2C and sideband signals on SFP+ connectors
    Port0_Tx_Fault                : in    std_logic;
    Port0_Tx_Disable              : out   std_logic;
    Port0_RS0                     : out   std_logic;
    Port0_RS1                     : out   std_logic;
    Port0_Mod_ABS                 : in    std_logic;
    Port0_SCL                     : inout std_logic;
    Port0_SDA                     : inout std_logic;
    Port0_Rx_LOS                  : in    std_logic;

    Port1_Tx_Fault                : in    std_logic;
    Port1_Tx_Disable              : out   std_logic;
    Port1_RS0                     : out   std_logic;
    Port1_RS1                     : out   std_logic;
    Port1_Mod_ABS                 : in    std_logic;
    Port1_SCL                     : inout std_logic;
    Port1_SDA                     : inout std_logic;
    Port1_Rx_LOS                  : in    std_logic;
    --vhook_nowarn Port*_S* Port*_RX_LOS Port*_Tx_Fault

    -- These are outputs that the CLIP asserts to drive the Active and Present LEDs
    -- on the SFP+ cage. Note these are active-high logic!
    LED_Port0Active               : out   std_logic;
    LED_Port1Active               : out   std_logic;
    LED_Port0Present              : out   std_logic;
    LED_Port1Present              : out   std_logic;

    -- 40 MHz Onboard Clock for use in the IO Socket
    -- For Aurora Cores generated in previous versions of Vivado, such as 2014.4,
    -- the Onboard Clock would have been sufficient to drive the init_clk. However,
    -- in Vivado 2015.4 init_clk must be driven with a minimum frequency of 50MHz.
    -- Thus, where SocketClk40 used to be implimented, DerivedClk50 is now used.
    SocketClk40                   : in    std_logic;
    --vhook_nowarn SocketClk40


    ----------------------------------------------------------------------------
    -- LVFPGA signals
    ----------------------------------------------------------------------------
    -- This is the collection of signals that appear in LabVIEW FPGA.
    --
    -- These signals are used to allow the user to interface with the CLIP
    -- from a high level perspective through LabVIEW as well as allowing the user
    -- to monitor the values associated with some of the internal signals
    --
    -- LabVIEW FPGA signals must use one of the following signal directions: {in, out}
    -- LabVIEW FPGA signals must use one of the following data types:
    --          std_logic
    --          std_logic_vector(7 downto 0)
    --          std_logic_vector(15 downto 0)
    --          std_logic_vector(31 downto 0)
    ----------------------------------------------------------------------------
    ------------------------ AXI Streaming TX Interface ------------------------
    -- The following signals are REQUIRED to be in the Port0UserClk domain:
    p0TxTData                     : in    std_logic_vector(63 downto 0);
    p0TxTValid                    : in    std_logic;
    p0TxTReady                    : out   std_logic;

    -- The following signals are REQUIRED to be in the Port1UserClk domain:
    p1TxTData                     : in    std_logic_vector(63 downto 0);
    p1TxTValid                    : in    std_logic;
    p1TxTReady                    : out   std_logic;

    ------------------------ AXI Streaming RX Interface ------------------------
    -- The following signals are REQUIRED to be in the Port0UserClk domain:
    p0RxTData                     : out   std_logic_vector(63 downto 0);
    p0RxTValid                    : out   std_logic;

    -- The following signals are REQUIRED to be in the Port1UserClk domain:
    p1RxTData                     : out   std_logic_vector(63 downto 0);
    p1RxTValid                    : out   std_logic;

    --------------------------- AXI4-Lite Interface ----------------------------
    -- This section is for MMCM and PLL Dynamic Reconfiguration(DRP) access

    -- AXI clk
    Lite_AXI_AClk                 : in    std_logic;

    -- This single AXI4-Lite Interface maps to two different endpoints.
    -- The address mapping values will be used in the
    -- Create AXI4-Lite Resources.vi in the LabVIEW FPGA diagram.
    -- Endpoint Address Width:     8
    -- Port0 GTXE2_CHANNEL Offset: 0
    -- Port1 GTXE2_CHANNEL Offset: 1

    -- The following signals are REQUIRED to be in the Lite_AXI_AClk domain:
    lManageAWAddr                 : in    std_logic_vector(31 downto 0);
    lManageAWValid                : in    std_logic;
    lManageAWReady                : out   std_logic;
    lManageWData                  : in    std_logic_vector(31 downto 0);
    lManageWValid                 : in    std_logic;
    lManageWReady                 : out   std_logic;
    lManageWStrb                  : in    std_logic_vector(3 downto 0);
    lManageBValid                 : out   std_logic;
    lManageBReady                 : in    std_logic;
    lManageBResp                  : out   std_logic_vector(1 downto 0);
    lManageARAddr                 : in    std_logic_vector(31 downto 0);
    lManageARValid                : in    std_logic;
    lManageARReady                : out   std_logic;
    lManageRData                  : out   std_logic_vector(31 downto 0);
    lManageRValid                 : out   std_logic;
    lManageRReady                 : in    std_logic;
    lManageRResp                  : out   std_logic_vector(1 downto 0);
    --vhook_nowarn lManageWStrb

    ----------------------------- Streaming Errors -----------------------------
    -- The following signals are REQUIRED to be in the Port0UserClk domain:
    p0HardError                   : out   std_logic;
    p0SoftError                   : out   std_logic;
    p0LaneUp                      : out   std_logic;
    p0ChannelUp                   : out   std_logic;

    -- The following signals are REQUIRED to be in the Port1UserClk domain:
    p1HardError                   : out   std_logic;
    p1SoftError                   : out   std_logic;
    p1LaneUp                      : out   std_logic;
    p1ChannelUp                   : out   std_logic;

    ---------------------------- Core Reset Status -----------------------------
    -- The following signal is REQUIRED to be in the Port0UserClk domain:
    p0SysResetOut                 : out   std_logic;

    -- The following signal is REQUIRED to be in the Port1UserClk domain:
    p1SysResetOut                 : out   std_logic;

    -- The following signals are REQUIRED to be in the DerivedClk50 Clock domain:
    dPort0LinkResetOut            : out   std_logic;
    dPort1LinkResetOut            : out   std_logic;

    ------------------------------ Signal Detect -------------------------------
    -- Detects signal from the high-speed serial connectors
    -- The following signal is REQUIRED to be in the Port0UserClk domain:
    p0SignalDetectPort0            : out   std_logic;

    -- The following signal is REQUIRED to be in the Port1UserClk domain:
    p1SignalDetectPort1            : out   std_logic;

    ----------------------------------- Misc -----------------------------------
    -- Asynchronous reset signal
    -- This signal *must* be present in the port interface for all IO Socket CLIPs.
    -- aReset should reset the CLIP logic whenever asserted high.
    -- It is assumed that this is signal that is not user-driven
    aReset                        : in    std_logic;

    -- AXI Streaming User Clock outputs (to LabVIEW FPGA diagram from I/O Socket)
    Port0UserClk                  : out   std_logic;
    Port1UserClk                  : out   std_logic;

    -- 50 MHz clock driven from LabVIEW, used instead of the Onboard Socket40 clock
    -- This specific CLIP expects a 50MHz clock to drive certain logic
    DerivedClk50                  : in    std_logic;

    -- Used to reset the Aurora cores post-powerup
    -- The following signals are REQUIRED to be in the DerivedClk50 domain:
    dPort0CoreReset               : in    std_logic;
    dPort1CoreReset               : in    std_logic

    );
end DualAuroraUsrpRio;


architecture rtl of DualAuroraUsrpRio is

  component IBUFDS_GTE2
    generic (
      CLKCM_CFG : boolean := TRUE;
      CLKRCV_TRST : boolean := TRUE;
      CLKSWING_CFG : bit_vector := "11");
    port (
      O : out std_logic;
      ODIV2 : out std_logic;
      CEB : in std_logic;
      I : in std_logic;
      IB : in std_logic);
  end component;
  --vhook_sigstart
  --vhook_sigend
  component OBUF
    port (
      I : in std_logic;
      O : out std_logic);
  end component;
  component ibuf
    port (
      I : in std_logic;
      O : out std_logic);
  end component;
  ---------------------------- Signal Declarations -----------------------------

  -- SLVs for the single lane port signals on the cores.
  signal Port0TxSlv_p, Port0TxSlv_n    : std_logic_vector(0 downto 0);
  signal Port0RxSlv_p, Port0RxSlv_n    : std_logic_vector(0 downto 0);
  signal p0LaneUpSlv                   : std_logic_vector(0 downto 0);
  signal Port1TxSlv_p, Port1TxSlv_n    : std_logic_vector(0 downto 0);
  signal Port1RxSlv_p, Port1RxSlv_n    : std_logic_vector(0 downto 0);
  signal p1LaneUpSlv                   : std_logic_vector(0 downto 0);

  -- Reversed range signals to accommodate the ports on the cores.
  signal p0RxTDataUp, p0TxTDataUp      : std_logic_vector(0 to 63) := (others =>'0');
  signal p1RxTDataUp, p1TxTDataUp      : std_logic_vector(0 to 63) := (others =>'0');

  -- Clock signals
  signal MGT_RefClk156p25MHz           : std_logic;
  signal Port0UserClkI, Port0TxOutClk, Port0_QPLL_RefInClk, Port0_QPLL_InClk,
         Port0SyncClk                  : std_logic;
  signal Port1UserClkI, Port1TxOutClk, Port1_QPLL_RefInClk, Port1_QPLL_InClk,
         Port1SyncClk                  : std_logic;
  --vhook_nowarn Port*_QPLL_InClk

  -- Internal Status and Control signals
  signal dPort0_QPLL_lock, dPort0_QPLL_RefClkLostIn, dPort0_MCMM_NotLocked,
         dPort0LinkResetOutI           : std_logic;
  signal p0SysResetOutI, p0SoftErr, p0HardErr,
         p0ChannelUpI                  : std_logic;
  signal aPort0_QPLL_ResetOut,
         aPort0_QPLL_LockIn            : std_logic;

  signal dPort1_QPLL_lock, dPort1_QPLL_RefClkLostIn, dPort1_MCMM_NotLocked,
         dPort1LinkResetOutI           : std_logic;
  signal p1SysResetOutI, p1SoftErr, p1HardErr,
         p1ChannelUpI                  : std_logic;
  signal aPort1_QPLL_ResetOut,
         aPort1_QPLL_LockIn            : std_logic;

  -- LED detect signals for front panel interfacing
  signal p0SignalDetectPort0Lcl        : std_logic;
  signal p1SignalDetectPort1Lcl        : std_logic;

  signal lLane_DRP_RdyOutSlv, lLane_DRP_EnInSlv,
         lLane_DRP_WeInSlv             : std_logic_vector(1 downto 0);

  -- AXI4-Lite Valid and Ready signal vectors
  signal lManageAWValidSlv, lManageAWReadySlv, lManageWValidSlv,
         lManageWReadySlv, lManageBValidSlv, lManageARValidSlv,
         lManageARReadySlv, lManageRValidSlv, lManageRReadySlv,
         lManageBReadySlv              : std_logic_vector(1 downto 0);

  -- Intermediate signals to allow user to read the output from the core
  signal p0RxTValidI, p0TxTReadyI      : std_logic;
  signal p1RxTValidI, p1TxTReadyI      : std_logic;

  -- RSD reset signals used to reset FSMs, logic, and counters
  signal adReset                       : std_logic;
  signal ap0Reset                      : std_logic;
  signal ap1Reset                      : std_logic;
  signal alReset                       : std_logic;
  signal alReset_n                     : std_logic;

  -- Intermediate signals between CoreResetFSM and their respective core
  signal dPort0CoreReset_pb,
         dPort0_PMA_Init               : std_logic;
  signal dPort1CoreReset_pb,
         dPort1_PMA_Init               : std_logic;

  -- AXI4-Lite Read Data vectors from the DRP endpoints in the cores
  subtype AxiData_t is std_logic_vector(31 downto 0);
  type AxiDataAry_t is array(natural range <>) of AxiData_t;
  signal lManageRDataLane                       : AxiDataAry_t(1 downto 0);
  signal lManageRDataLcl                        : AxiData_t;

  -- MGT Lane DRP signals
  subtype DrpAddr_t is std_logic_vector(8 downto 0);
  type DrpAddrAry_t is array(natural range <>) of DrpAddr_t;
  signal lLane_DRP_AddrIn                       : DrpAddrAry_t(1 downto 0);

  subtype DrpData_t is std_logic_vector(15 downto 0);
  type DrpDataAry_t is array(natural range <>) of DrpData_t;
  signal lLane_DRPDI_In, lLane_DRPDO_Out        : DrpDataAry_t(1 downto 0);


  --------------------------- Component Declarations ---------------------------
  component AuroraCore64b66b
    port (
      rxp             : in    std_logic_vector(0 downto 0);
      rxn             : in    std_logic_vector(0 downto 0);
      refclk1_in      : in    std_logic;
      user_clk        : in    std_logic;
      sync_clk        : in    std_logic;
      power_down      : in    std_logic;
      pma_init        : in    std_logic;
      loopback        : in    std_logic_vector(2 downto 0);
      txp             : out   std_logic_vector(0 downto 0);
      txn             : out   std_logic_vector(0 downto 0);
      hard_err        : out   std_logic;
      soft_err        : out   std_logic;
      channel_up      : out   std_logic;
      lane_up         : out   std_logic_vector(0 downto 0);
      tx_out_clk      : out   std_logic;
      drp_clk_in      : in    std_logic;
      gt_pll_lock     : out   std_logic;
      s_axi_tx_tdata  : in    std_logic_vector(0 to 63);
      s_axi_tx_tvalid : in    std_logic;
      s_axi_tx_tready : out   std_logic;
      m_axi_rx_tdata  : out   std_logic_vector(0 to 63);
      m_axi_rx_tvalid : out   std_logic;
      mmcm_not_locked : in    std_logic;
      drpaddr_in      : in    std_logic_vector(8 downto 0);
      drpdi_in        : in    std_logic_vector(15 downto 0);
      qpll_drpaddr_in : in    std_logic_vector(7 downto 0);
      qpll_drpdi_in   : in    std_logic_vector(15 downto 0);
      drprdy_out      : out   std_logic;
      drpen_in        : in    std_logic;
      drpwe_in        : in    std_logic;
      qpll_drprdy_out : out   std_logic;
      qpll_drpen_in   : in    std_logic;
      qpll_drpwe_in   : in    std_logic;
      drpdo_out       : out   std_logic_vector(15 downto 0);
      qpll_drpdo_out  : out   std_logic_vector(15 downto 0);
      init_clk        : in    std_logic;
      link_reset_out  : out   std_logic;
      gt_qpllclk_quad1_in        : in    std_logic;
      gt_qpllrefclk_quad1_in     : in    std_logic;
      gt_to_common_qpllreset_out : out   std_logic;
      gt_qplllock_in             : in    std_logic;
      gt_qpllrefclklost_in       : in    std_logic;
      gt_rxcdrovrden_in          : in    std_logic;
      sys_reset_out   : out   std_logic;
      reset_pb        : in    std_logic
    );
  end component;
  attribute syn_black_box                      : boolean;
  attribute syn_black_box of AuroraCore64b66b  : component is true;

  component AuroraCore64b66b_gt_common_wrapper
    port (
      gt_qpllclk_quad1_out    : out   std_logic;
      gt_qpllrefclk_quad1_out : out   std_logic;
      gt0_gtrefclk0_common_in : in    std_logic;
      gt0_qplllock_out        : out   std_logic;
      gt0_qpllreset_in        : in    std_logic;
      gt0_qplllockdetclk_in   : in    std_logic;
      gt0_qpllrefclklost_out  : out   std_logic
    );
  end component;
  attribute syn_black_box of AuroraCore64b66b_gt_common_wrapper   : component is true;

  component AuroraCore64b66b_CLOCK_MODULE
    port (
      init_clk_p              : in    std_logic;
      init_clk_n              : in    std_logic;
      init_clk_o              : out   std_logic;
      clk                     : in    std_logic;
      clk_locked              : in    std_logic;
      user_clk                : out   std_logic;
      sync_clk                : out   std_logic;
      mmcm_not_locked         : out   std_logic
    );
  end component;
  attribute syn_black_box of AuroraCore64b66b_CLOCK_MODULE        : component is true;

  component OBUFDS
    port (
      O               : out   std_logic;
      OB              : out   std_logic;
      I               : in    std_logic);
  end component;

  component ResetSyncDeassertion
    port (
      aReset          : in    std_logic;
      Clk             : in    std_logic;
      acReset         : out   std_logic);
  end component;

  --------------------------------- Functions ----------------------------------
  -- The following function reverses the bits of the input and returns it
  function reverse (arg : std_logic_vector) return std_logic_vector is
    variable RetVal : std_logic_vector(arg'reverse_range) := (others => '0');

  begin
      for index in arg'range loop
        RetVal(index) := arg(index);
      end loop;
    return RetVal;
  end reverse;


begin

  ---------------------------------------------------------------------------------------
  -- Transmit (Output) Buffers
  ---------------------------------------------------------------------------------------
  Port0TxBuf_p : OBUF
    port map (
      I => Port0TxSlv_p(0),           -- in  std_logic
      O => Port0_TX_p);               -- out std_logic

  Port0TxBuf_n : OBUF
    port map (
      I => Port0TxSlv_n(0),           -- in  std_logic
      O => Port0_TX_n);               -- out std_logic

  Port1TxBuf_p : OBUF
    port map (
      I => Port1TxSlv_p(0),           -- in  std_logic
      O => Port1_TX_p);               -- out std_logic

  Port1TxBuf_n : OBUF
    port map (
      I => Port1TxSlv_n(0),           -- in  std_logic
      O => Port1_TX_n);               -- out std_logic

  ---------------------------------------------------------------------------------------
  -- Receive (Input) Buffers
  ---------------------------------------------------------------------------------------
  Port0RxBuf_p : ibuf
    port map (
      I => Port0_RX_p,                -- in  std_logic
      O => Port0RxSlv_p(0));          -- out std_logi

  Port0RxBuf_n : ibuf
    port map (
      I => Port0_RX_n,                -- in  std_logic
      O => Port0RxSlv_n(0));          -- out std_logic

  Port1RxBuf_p : ibuf
    port map (
      I => Port1_RX_p,                -- in  std_logic
      O => Port1RxSlv_p(0));          -- out std_logic

  Port1RxBuf_n : ibuf
    port map (
      I => Port1_RX_n,                -- in  std_logic
      O => Port1RxSlv_n(0));          -- out std_logic


  -- Interfacing the transceiver pins with signals used by the core
  -- Port0_TX_p       <= Port0TxSlv_p(0);
  -- Port0_TX_n       <= Port0TxSlv_n(0);
  -- Port1_TX_p       <= Port1TxSlv_p(0);
  -- Port1_TX_n       <= Port1TxSlv_n(0);

  -- Port0RxSlv_p(0)  <= Port0_RX_p;
  -- Port0RxSlv_n(0)  <= Port0_RX_n;
  -- Port1RxSlv_p(0)  <= Port1_RX_p;
  -- Port1RxSlv_n(0)  <= Port1_RX_n;

  -- Rate Select: RS0 and RS1 are always set to 1 for operation above 4.25 Gbps
  -- We are operating at 10.3125 Gbps
  Port0_RS0        <= '1';
  Port1_RS0        <= '1';
  Port0_RS1        <= '1';
  Port1_RS1        <= '1';

  -- Enabling Tx for both ports
  Port1_Tx_Disable <= '0';
  Port0_Tx_Disable <= '0';

  -- Routing local signals to the top-level
  p0RxTValid       <= p0RxTValidI;
  p0TxTReady       <= p0TxTReadyI;
  p1RxTValid       <= p1RxTValidI;
  p1TxTReady       <= p1TxTReadyI;


  ------------------------------------------------------------------------------
  -- Clock Domain Crossing - RSD Resets
  ------------------------------------------------------------------------------
  --
  -- The following block contains the logic used to to ensure proper handling
  -- for asynchronous resets with synchronous de-assertion.
  --
  ------------------------------------------------------------------------------
  -- RSD reset for DerivedClk50 clock domain
  RSD_Derived50Clk : ResetSyncDeassertion
  port map(
      aReset  => aReset,
      Clk     => DerivedClk50,
      acReset => adReset
      );

  -- RSD reset for Port0UserClk clock domain
  RSD_Port0Clk     : ResetSyncDeassertion
  port map(
      aReset  => aReset,
      Clk     => Port0UserClkI,
      acReset => ap0Reset
      );

  -- RSD reset for Port1UserClk clock domain
  RSD_Port1Clk     : ResetSyncDeassertion
  port map(
      aReset  => aReset,
      Clk     => Port1UserClkI,
      acReset => ap1Reset
      );

  -- RSD reset for Lite_AXI_AClk clock domain
  RSD_Lite_AXI_Clk : ResetSyncDeassertion
  port map(
      aReset  => aReset,
      Clk     => Lite_AXI_AClk,
      acReset => alReset
      );

  -- Since the Lite_AXI_AClk reset is active low, invert it
  alReset_n   <= (not alReset);


  ------------------------------------------------------------------------------
  -- Clock Domain Crossing - LEDs
  ------------------------------------------------------------------------------
  -- There were no explicit instructions on how to drive the LEDs using a signal
  -- detect from the Aurora Core Product User Guide. However, in the Xilinx
  -- documentation for the PCS/PMA core (PG068), it recommends driving signal_detect
  -- with the NOR of MODDEF0 (ModAbs = Module Absent) and LOS (loss of signal).
  -- Since we also use this signal to drive LEDs and Window ports, we first
  -- synchronize all inputs to the common clock and reset.
  --
  -- Although the implementation of the signal detect was not specifically stated
  -- for the Aurora Core, the code uses the same concept as the
  -- PCS/PMA core. The theory was tested, and proven to work.
  --
  -- SFP+ Low Speed signals per SFF-8431 specification.
  ------------------------------------------------------------------------------
  ---------------- LED Signal Port 0 User Clock Domain Crossing ----------------
  SyncPort0RegBlock: block
    signal p0Port0ModAbs      : std_logic;
    signal p0Port0ModAbs_ms   : std_logic;
    signal p0Port0RxLos       : std_logic;
    signal p0Port0RxLos_ms    : std_logic;

    attribute ASYNC_REG : string;
    attribute ASYNC_REG of p0Port0ModAbs          : signal is "true";
    attribute ASYNC_REG of p0Port0ModAbs_ms       : signal is "true";
    attribute ASYNC_REG of p0Port0RxLos           : signal is "true";
    attribute ASYNC_REG of p0Port0RxLos_ms        : signal is "true";

    -- Keeps the synthesizer from optimizing into a shift register.
    attribute SHREG_EXTRACT : string;
    attribute SHREG_EXTRACT of p0Port0ModAbs      : signal is "no";
    attribute SHREG_EXTRACT of p0Port0ModAbs_ms   : signal is "no";
    attribute SHREG_EXTRACT of p0Port0RxLos       : signal is "no";
    attribute SHREG_EXTRACT of p0Port0RxLos_ms    : signal is "no";
  begin
    SyncReg0: process(ap0Reset, Port0UserClkI)
    begin
      if (ap0Reset = '1') then
        -- ModAbs and RxLos both reset to '1', meaning the module starts by assuming
        -- the module is absent and there is no signal present.
        p0Port0ModAbs_ms       <= '1';
        p0Port0ModAbs          <= '1';
        p0Port0RxLos_ms        <= '1';
        p0Port0RxLos           <= '1';

        -- Based on the above reset values, the signal detect value will be false after
        -- coming out of reset.
        p0SignalDetectPort0Lcl <= '0';

        -- Add another flop stage to reliably place false path constraints on this flop.
        -- The signal is driven to the top-level LabVIEW interface
        p0SignalDetectPort0    <= '0';

      elsif rising_edge(Port0UserClkI) then
        p0Port0ModAbs_ms       <= Port0_Mod_ABS;
        p0Port0ModAbs          <= p0Port0ModAbs_ms;

        p0Port0RxLos_ms        <= Port0_Rx_LOS;
        p0Port0RxLos           <= p0Port0RxLos_ms;

        p0SignalDetectPort0Lcl <= p0Port0ModAbs nor p0Port0RxLos;

        -- Send signal detect to LabVIEW.
        p0SignalDetectPort0    <= p0SignalDetectPort0Lcl;
      end if;
    end process SyncReg0;

  end block SyncPort0RegBlock;

  ---------------- LED Signal Port 1 User Clock Domain Crossing ----------------
  SyncPort1RegBlock: block
    signal p1Port1ModAbs     : std_logic;
    signal p1Port1ModAbs_ms  : std_logic;
    signal p1Port1RxLos      : std_logic;
    signal p1Port1RxLos_ms   : std_logic;

    -- In this application, ASYNC_REG is used to specify that the following registers
    -- are a synchronizing register within a synchronization chain.
    attribute ASYNC_REG : string;
    attribute ASYNC_REG of p1Port1ModAbs        : signal is "true";
    attribute ASYNC_REG of p1Port1ModAbs_ms     : signal is "true";
    attribute ASYNC_REG of p1Port1RxLos         : signal is "true";
    attribute ASYNC_REG of p1Port1RxLos_ms      : signal is "true";

    -- Keeps the synthesizer from optimizing into a shift register.
    attribute SHREG_EXTRACT : string;
    attribute SHREG_EXTRACT of p1Port1ModAbs    : signal is "no";
    attribute SHREG_EXTRACT of p1Port1ModAbs_ms : signal is "no";
    attribute SHREG_EXTRACT of p1Port1RxLos     : signal is "no";
    attribute SHREG_EXTRACT of p1Port1RxLos_ms  : signal is "no";
  begin
    SyncReg1: process(ap1Reset, Port1UserClkI)
    begin
      if (ap1Reset = '1') then
        -- ModAbs and RxLos both reset to '1', meaning the module starts by assuming
        -- the module is absent and there is no signal present.
        p1Port1ModAbs_ms       <= '1';
        p1Port1ModAbs          <= '1';
        p1Port1RxLos_ms        <= '1';
        p1Port1RxLos           <= '1';

        -- Based on the above reset values, the signal detect value will be false after
        -- coming out of reset.
        p1SignalDetectPort1Lcl <= '0';

        -- Add another flop stage to reliably place false path constraints on this flop.
        -- The signal is driven to the top-level LabVIEW interface
        p1SignalDetectPort1    <= '0';

      elsif rising_edge(Port1UserClkI) then
        p1Port1ModAbs_ms       <= Port1_Mod_ABS;
        p1Port1ModAbs          <= p1Port1ModAbs_ms;

        p1Port1RxLos_ms        <= Port1_Rx_LOS;
        p1Port1RxLos           <= p1Port1RxLos_ms;

        p1SignalDetectPort1Lcl <= p1Port1ModAbs nor p1Port1RxLos;

        -- Send signal detect to LabVIEW.
        p1SignalDetectPort1    <= p1SignalDetectPort1Lcl;
      end if;
    end process SyncReg1;

  end block SyncPort1RegBlock;


  ------------------------------------------------------------------------------
  -- User Interface - CLIP Reset Signals
  ------------------------------------------------------------------------------
  ClipResetOut : process (adReset, DerivedClk50) is
  begin
    if (adReset = '1') then
      dPort0LinkResetOut <= '1';
      dPort1LinkResetOut <= '1';
    elsif rising_edge(DerivedClk50) then
      dPort0LinkResetOut <= dPort0LinkResetOutI;
      dPort1LinkResetOut <= dPort1LinkResetOutI;
    end if;
  end process ClipResetOut;


  ------------------------------------------------------------------------------
  -- Core Reset Sequence
  ------------------------------------------------------------------------------
  --
  -- The following are declarations of the CoreResetFSM component which is
  -- used for the reset logic of the Aurora 64B/66B. It will be used to ensure
  -- proper resetting in accordance with the Xilinx Product User Guide (PG074) v11.1
  -- page 61.
  ------------------------------------------------------------------------------
  -- Reset Sequence for Core 0
  --vhook_e CoreResetFSM Port0CoreResetFSM
  --vhook_g k*  open
  --vhook_a dCoreUserReset dPort0CoreReset
  --vhook_a dPmaInit       dPort0_PMA_Init
  --vhook_a dResetPb       dPort0CoreReset_pb
  --vhook_a dCounterDbg    open
  Port0CoreResetFSM: entity work.CoreResetFSM (rtl)
    generic map (
      kCounterWidth             => open,  -- in  positive := 26
      kClksBtwResetsDeassertion => open,  -- in  positive range 1 to 1023 := 4
      kClksBtwResetsAssertion   => open)  -- in  positive range 1 to 1023 := 40
    port map (
      adReset        => adReset,             -- in  std_logic
      DerivedClk50   => DerivedClk50,        -- in  std_logic
      dCoreUserReset => dPort0CoreReset,     -- in  std_logic
      dPmaInit       => dPort0_PMA_Init,     -- out std_logic
      dResetPb       => dPort0CoreReset_pb,  -- out std_logic
      dCounterDbg    => open);               -- out unsigned((kCounterWidth-1)downto 0)

  -- Reset Sequence for Core 1
  --vhook_e CoreResetFSM Port1CoreResetFSM
  --vhook_g k*  open
  --vhook_a dCoreUserReset dPort1CoreReset
  --vhook_a dPmaInit       dPort1_PMA_Init
  --vhook_a dResetPb       dPort1CoreReset_pb
  --vhook_a dCounterDbg    open
  Port1CoreResetFSM: entity work.CoreResetFSM (rtl)
    generic map (
      kCounterWidth             => open,  -- in  positive := 26
      kClksBtwResetsDeassertion => open,  -- in  positive range 1 to 1023 := 4
      kClksBtwResetsAssertion   => open)  -- in  positive range 1 to 1023 := 40
    port map (
      adReset        => adReset,             -- in  std_logic
      DerivedClk50   => DerivedClk50,        -- in  std_logic
      dCoreUserReset => dPort1CoreReset,     -- in  std_logic
      dPmaInit       => dPort1_PMA_Init,     -- out std_logic
      dResetPb       => dPort1CoreReset_pb,  -- out std_logic
      dCounterDbg    => open);               -- out unsigned((kCounterWidth-1)downto 0)


  ------------------------------------------------------------------------------
  -- LED Control Sequence
  ------------------------------------------------------------------------------
  --
  -- The following block contains the logic for driving the external LEDs - Signal
  -- Present, and Signal Active - for both Port 0 and Port 1
  --
  -- !!! SAFE STATE MACHINE AND COUNTER STARTUP !!!
  -- The following state machines and counters have a safe startup because they
  -- are driven by an RSD reset.
  --
  ------------------------------------------------------------------------------
  LedsBlock : block
    signal p0Port0ActiveLed : std_logic;
    signal p1Port1ActiveLed : std_logic;

    -- Each clock tick is 161.1328125 MHz ~= 6.2 ns, so we require
    -- log2(50 ms/6.2 ns) ~= 23 bits to meet the roughly 50 ms flashing period.
    signal p0Port0LedCount,
           p1Port1LedCount  : unsigned(22 downto 0);

    type   LedState_t is (Idle, Accessed, WaitForStart, WaitForEnd);
    signal p0Port0LedState  : LedState_t;
    signal p1Port1LedState  : LedState_t;

  begin
    --------------------------- LED Port 0 FSM ---------------------------------
    -- If a SFP+ cable is connected, set the Port 0 Present LEDs.
    -- If there is activity on the cable, set the Port 0 Active LEDs.
    LedRegPort0: process(ap0Reset, Port0UserClkI)
    begin

      if (ap0Reset = '1') then
        p0Port0ActiveLed  <= '0';
        p0Port0LedCount   <= (others => '0');
        p0Port0LedState   <= Idle;

      elsif rising_edge(Port0UserClkI) then

        -- Keep the Active LED on for at least 50-150ms so it is visible to the user.
        -- Set up a port specific counter that starts running when the specified port's
        -- cable is present. This is an easy way to guarantee safe startup, and that
        -- the active LED will never assert if the present LED is not asserted.

        if (p0SignalDetectPort0Lcl = '1') then
          -- Counter will continue to count and roll over as Port 0's cable is present.
          p0Port0LedCount    <= p0Port0LedCount + 1;
        end if;

        -- Default state is the LED turned on, although since it starts in Idle the
        -- LED is turned off until the FSM transitions out of Idle.
        p0Port0ActiveLed     <= '1';

        case p0Port0LedState is
          when Idle =>
            -- Any other state allows the default statement above
            -- to take control and turn on the LED.
            p0Port0ActiveLed <= '0';

            -- Determine if the links are active: when we receive data or when we are
            -- actively transmitting data.
            if ((p0RxTValidI = '1') or
               (p0TxTValid   = '1' and p0TxTReadyI = '1')) and
               (p0SignalDetectPort0Lcl = '1') then
              p0Port0LedState <= Accessed;
            end if;

          when Accessed =>

            if (p0Port0LedCount(p0Port0LedCount'high) = '0') then
              p0Port0LedState <= WaitForStart;
            end if;

          when WaitForStart =>

            if (p0Port0LedCount(p0Port0LedCount'high) = '1') then
              p0Port0LedState <= WaitForEnd;
            end if;

          when WaitForEnd =>

            if (p0Port0LedCount(p0Port0LedCount'high) = '0') then
              p0Port0LedState <= Idle;
            end if;

          -- Default state
          when others =>
            p0Port0LedState   <= Idle;
          end case;

        end if;
      end process LedRegPort0;


      ----------------------------- LED Port 1 FSM -----------------------------
      -- If a SFP+ cable is connected, set the Port 1 Present LEDs.
      -- If there is activity on the cable, set the Port 1 Active LEDs.
      LedRegPort1: process(ap1Reset, Port1UserClkI)
      begin

        if (ap1Reset = '1') then
          p1Port1ActiveLed  <= '0';
          p1Port1LedCount   <= (others => '0');
          p1Port1LedState   <= Idle;

        elsif rising_edge(Port1UserClkI) then

          -- Keep the Active LED on for at least 50-150ms so it is visible to the user.
          -- Set up a port specific counter that starts running when the specified port's
          -- cable is present. This is an easy way to guarantee safe startup, and that
          -- the active LED will never assert if the present LED is not asserted.

          if (p1SignalDetectPort1Lcl = '1') then
            -- Counter will continue to count and roll over as Port 1's cable is present.
            p1Port1LedCount <= p1Port1LedCount + 1;
          end if;

          -- Default state is the LED turned on, although since it starts in Idle the
          -- LED is turned off until the FSM transitions out of Idle.
          p1Port1ActiveLed   <= '1';

        case p1Port1LedState is
          when Idle =>
            -- Any other state allows the default statement above
            -- to take control and turn on the LED.
            p1Port1ActiveLed <= '0';

            -- Determine if the links are active: when we receive data or when we are
            -- actively transmitting data.
            if ((p1RxTValidI = '1') or
               (p1TxTValid   = '1' and p1TxTReadyI = '1')) and
               (p1SignalDetectPort1Lcl = '1') then
              p1Port1LedState <= Accessed;
            end if;

          -- The following three states are used for the blinking mechanics
          when Accessed =>

            if (p1Port1LedCount(p1Port1LedCount'high) = '0') then
              p1Port1LedState <= WaitForStart;
            end if;

          when WaitForStart =>

            if (p1Port1LedCount(p1Port1LedCount'high) = '1') then
              p1Port1LedState <= WaitForEnd;
            end if;

          when WaitForEnd =>

            if (p1Port1LedCount(p1Port1LedCount'high) = '0') then
              p1Port1LedState <= Idle;
            end if;

          when others =>
            p1Port1LedState   <= Idle;
        end case;

      end if;
    end process LedRegPort1;

    -- Locals to outputs.
    LED_Port0Active  <= p0Port0ActiveLed;
    LED_Port1Active  <= p1Port1ActiveLed;

    -- When signal is detected on the cable, a cable should be present, so we illuminate
    -- the present LED.
    LED_Port0Present <= p0SignalDetectPort0Lcl;
    LED_Port1Present <= p1SignalDetectPort1Lcl;

  end block;


  ------------------------------------------------------------------------------
  -- AuroraBlock
  ------------------------------------------------------------------------------
  AuroraBlock : block
  begin

    -- Routing local signals to the top-level - LabVIEW
    -- This enables the user to implement their design in the proper clock domain
    Port0UserClk <= Port0UserClkI;
    Port1UserClk <= Port1UserClkI;

    ----------------------------------------------------------------------------
    -- Register User I/O
    ----------------------------------------------------------------------------
    -- Register outputs driven from the core to LabVIEW for user debug convenience
    Port0RegUserOutputs : process(ap0Reset, Port0UserClkI)
    begin
      if (ap0Reset = '1') then
        p0HardError      <= '0';
        p0SoftError      <= '0';
        p0LaneUp         <= '0';
        p0ChannelUp      <= '0';
        p0SysResetOut    <= '1';
      elsif rising_edge(Port0UserClkI) then
        p0HardError      <= p0HardErr;
        p0SoftError      <= p0SoftErr;
        p0LaneUp         <= p0LaneUpSlv(0);
        p0ChannelUp      <= p0ChannelUpI;
        p0SysResetOut    <= p0SysResetOutI;
      end if;
    end process Port0RegUserOutputs;

    Port1RegUserOutputs : process(ap1Reset, Port1UserClkI)
    begin
      if (ap1Reset = '1') then
        p1HardError      <= '0';
        p1SoftError      <= '0';
        p1LaneUp         <= '0';
        p1ChannelUp      <= '0';
        p1SysResetOut    <= '1';
      elsif rising_edge(Port1UserClkI) then
        p1HardError      <= p1HardErr;
        p1SoftError      <= p1SoftErr;
        p1LaneUp         <= p1LaneUpSlv(0);
        p1ChannelUp      <= p1ChannelUpI;
        p1SysResetOut    <= p1SysResetOutI;
      end if;
    end process Port1RegUserOutputs;


    ----------------------------------------------------------------------------
    -- AXI4-Lite and DRP Handlers
    ----------------------------------------------------------------------------
    -------------------------- AXI4_Lite Address Map ---------------------------
    -- This component uses a single AXI4-Lite bus to index into multiple
    -- AXI4-Lite slaves. It uses the kNumEndpoints generic to determine the size
    -- of the select vector and the size of the slave vectors. The kAddrSelectLsb
    -- generic is used to determine the offset into the AXI4-Lite address vector
    -- for the selection vector. The select value is updated whenever read or
    -- write address valid is strobed with the priority going to read address valid.
    -- This component does not route read or write data through it.
    ----------------------------------------------------------------------------
    AXI4_LiteAddressMap : entity work.USRP_RIO_AXI4_Lite_Address_Map(rtl)
      generic map (
        kNumEndpoints  => 2,
        kAddrSelectLsb => 9
      )
      port map (
        s_aclk              => Lite_AXI_AClk,
        aReset_n            => alReset_n,
        s_axi_awaddr        => lManageAWAddr,
        s_axi_awvalid       => lManageAWValid,
        s_axi_awready       => lManageAWReady,
        s_axi_wvalid        => lManageWValid,
        s_axi_wready        => lManageWReady,
        s_axi_bvalid        => lManageBValid,
        s_axi_bready        => lManageBReady,
        s_axi_araddr        => lManageARAddr,
        s_axi_arvalid       => lManageARValid,
        s_axi_arready       => lManageARReady,
        s_axi_rdata         => lManageRData,
        s_axi_rvalid        => lManageRValid,
        s_axi_rready        => lManageRReady,
        s_axi_awvalid_slv   => lManageAWValidSlv,
        s_axi_awready_slv   => lManageAWReadySlv,
        s_axi_wvalid_slv    => lManageWValidSlv,
        s_axi_wready_slv    => lManageWReadySlv,
        s_axi_bvalid_slv    => lManageBValidSlv,
        s_axi_bready_slv    => lManageBReadySlv,
        s_axi_arvalid_slv   => lManageARValidSlv,
        s_axi_arready_slv   => lManageARReadySlv,
        s_axi_rdata_in      => lManageRDataLcl,
        s_axi_rvalid_slv    => lManageRValidSlv,
        s_axi_rready_slv    => lManageRReadySlv
      );

    ---------------------------- AXI4_Lite To DRP ----------------------------
    -- This component does a simple translation from the AXI4-Lite bus to the
    -- Xilinx DRP bus. It has two simple state machines for read and write
    -- transactions to guarantee compatibility with the AXI4-Lite and DRP protocols.
    --------------------------------------------------------------------------
    GenAxiDrplanes : for i in 0 to 1 generate
      Port0Lane_AXI4_LiteToDRP : entity work.USRP_RIO_AXI4_Lite_to_DRP(rtl)
        port map (
          s_aclk            => Lite_AXI_AClk,
          aReset_n          => alReset_n,
          s_axi_awaddr      => lManageAWAddr,
          s_axi_awvalid     => lManageAWValidSlv(i),
          s_axi_awready     => lManageAWReadySlv(i),
          s_axi_wdata       => lManageWData,
          s_axi_wvalid      => lManageWValidSlv(i),
          s_axi_wready      => lManageWReadySlv(i),
          s_axi_bready      => lManageBReadySlv(i),
          s_axi_bvalid      => lManageBValidSlv(i),
          s_axi_araddr      => lManageARAddr,
          s_axi_arvalid     => lManageARValidSlv(i),
          s_axi_arready     => lManageARReadySlv(i),
          s_axi_rdata       => lManageRDataLane(i),
          s_axi_rready      => lManageRReadySlv(i),
          s_axi_rvalid      => lManageRValidSlv(i),
          drpaddr_in        => lLane_DRP_AddrIn(i),
          drpdi_in          => lLane_DRPDI_In(i),
          drpdo_out         => lLane_DRPDO_Out(i),
          drprdy_out        => lLane_DRP_RdyOutSlv(i),
          drpen_in          => lLane_DRP_EnInSlv(i),
          drpwe_in          => lLane_DRP_WeInSlv(i)
        );
    end generate;

    lManageRResp    <= "00";
    lManageBResp    <= "00";
    lManageRDataLcl <= lManageRDataLane(1) or lManageRDataLane(0);


    ----------------------------------------------------------------------------
    -- Module Instantiations
    ----------------------------------------------------------------------------
    ----------------------------- Shared Modules -------------------------------
    -- Dedicated MGT Input Clock Buffer
    MGT_RefClk156p25MHzIBuf : IBUFDS_GTE2
      port map (
        O                          => MGT_RefClk156p25MHz,
        ODIV2                      => open,
        CEB                        => '0',
        I                          => MGT_RefClk156p25MHz_p,
        IB                         => MGT_RefClk156p25MHz_n
      );

    ------------------------------ Port0 Modules -------------------------------
    -- Instantiates the QPLL wrapper
    Port0CommonWrapper : AuroraCore64b66b_gt_common_wrapper
      port map (
        gt_qpllclk_quad1_out       => Port0_QPLL_InClk,
        gt_qpllrefclk_quad1_out    => Port0_QPLL_RefInClk,
        gt0_gtrefclk0_common_in    => MGT_RefClk156p25MHz,
        gt0_qplllock_out           => aPort0_QPLL_LockIn,
        gt0_qpllreset_in           => aPort0_QPLL_ResetOut,
        gt0_qplllockdetclk_in      => DerivedClk50,
        gt0_qpllrefclklost_out     => dPort0_QPLL_RefClkLostIn
      );

    -- Instantiate a clock module for clock division.
    Port0ClockModule : AuroraCore64b66b_CLOCK_MODULE
      port map (
        init_clk_p                 => '0',
        init_clk_n                 => '0',
        init_clk_o                 => open,
        clk                        => Port0TxOutClk,
        clk_locked                 => dPort0_QPLL_lock,
        user_clk                   => Port0UserClkI,
        sync_clk                   => Port0SyncClk,
        mmcm_not_locked            => dPort0_MCMM_NotLocked
      );

    -- Instantiate the Aurora 64b66b Core
    Port0AuroraCore64b66b : AuroraCore64b66b
      port map (
        rxp                        => Port0RxSlv_p,
        rxn                        => Port0RxSlv_n,
        refclk1_in                 => MGT_RefClk156p25MHz,
        user_clk                   => Port0UserClkI,
        sync_clk                   => Port0SyncClk,
        power_down                 => '0',
        pma_init                   => dPort0_PMA_Init,
        loopback                   => (others => '0'),
        txp                        => Port0TxSlv_p,
        txn                        => Port0TxSlv_n,
        hard_err                   => p0HardErr,
        soft_err                   => p0SoftErr,
        channel_up                 => p0ChannelUpI,
        lane_up                    => p0LaneUpSlv,
        tx_out_clk                 => Port0TxOutClk,
        drp_clk_in                 => Lite_AXI_AClk,
        gt_pll_lock                => dPort0_QPLL_lock,
        s_axi_tx_tdata             => p0TxTDataUp,
        s_axi_tx_tvalid            => p0TxTValid,
        s_axi_tx_tready            => p0TxTReadyI,
        m_axi_rx_tdata             => p0RxTDataUp,
        m_axi_rx_tvalid            => p0RxTValidI,
        mmcm_not_locked            => dPort0_MCMM_NotLocked,
        drpaddr_in                 => lLane_DRP_AddrIn(0),
        drpdi_in                   => lLane_DRPDI_In(0),
        qpll_drpaddr_in            => (others => '0'),
        qpll_drpdi_in              => (others => '0'),
        drprdy_out                 => lLane_DRP_RdyOutSlv(0),
        drpen_in                   => lLane_DRP_EnInSlv(0),
        drpwe_in                   => lLane_DRP_WeInSlv(0),
        qpll_drprdy_out            => open,
        qpll_drpen_in              => '0',
        qpll_drpwe_in              => '0',
        drpdo_out                  => lLane_DRPDO_Out(0),
        qpll_drpdo_out             => open,
        init_clk                   => DerivedClk50,
        link_reset_out             => dPort0LinkResetOutI,
        gt_qpllclk_quad1_in        => Port0_QPLL_InClk,
        gt_qpllrefclk_quad1_in     => Port0_QPLL_RefInClk,
        gt_to_common_qpllreset_out => aPort0_QPLL_ResetOut,
        gt_qplllock_in             => aPort0_QPLL_LockIn,
        gt_qpllrefclklost_in       => dPort0_QPLL_RefClkLostIn,
        gt_rxcdrovrden_in          => '0',
        sys_reset_out              => p0SysResetOutI,
        reset_pb                   => dPort0CoreReset_pb
      );

    -- Reversing the Data Values
    -- To transmit data, the Lsb is left-most
    p0TxTDataUp <= reverse(p0TxTData);
    p0RxTData   <= reverse(p0RxTDataUp);


    ------------------------------ Port0 Modules -------------------------------
    -- Instantiate the QPLL wrapper.
    Port1CommonWrapper : AuroraCore64b66b_gt_common_wrapper
      port map (
        gt_qpllclk_quad1_out       => Port1_QPLL_InClk,
        gt_qpllrefclk_quad1_out    => Port1_QPLL_RefInClk,
        gt0_gtrefclk0_common_in    => MGT_RefClk156p25MHz,
        gt0_qplllock_out           => aPort1_QPLL_LockIn,
        gt0_qpllreset_in           => aPort1_QPLL_ResetOut,
        gt0_qplllockdetclk_in      => DerivedClk50,
        gt0_qpllrefclklost_out     => dPort1_QPLL_RefClkLostIn
      );

    -- Instantiate a clock module for clock division.
    Port1ClockModule : AuroraCore64b66b_CLOCK_MODULE
      port map (
        init_clk_p                 => '0',
        init_clk_n                 => '0',
        init_clk_o                 => open,
        clk                        => Port1TxOutClk,
        clk_locked                 => dPort1_QPLL_lock,
        user_clk                   => Port1UserClkI,
        sync_clk                   => Port1SyncClk,
        mmcm_not_locked            => dPort1_MCMM_NotLocked
      );

    -- Instantiate the Aurora 64b66b Core
    Port1AuroraCore64b66b : AuroraCore64b66b
      port map (
        rxp                        => Port1RxSlv_p,
        rxn                        => Port1RxSlv_n,
        refclk1_in                 => MGT_RefClk156p25MHz,
        user_clk                   => Port1UserClkI,
        sync_clk                   => Port1SyncClk,
        power_down                 => '0',
        pma_init                   => dPort1_PMA_Init,
        loopback                   => (others => '0'),
        txp                        => Port1TxSlv_p,
        txn                        => Port1TxSlv_n,
        hard_err                   => p1HardErr,
        soft_err                   => p1SoftErr,
        channel_up                 => p1ChannelUpI,
        lane_up                    => p1LaneUpSlv,
        tx_out_clk                 => Port1TxOutClk,
        drp_clk_in                 => Lite_AXI_AClk,
        gt_pll_lock                => dPort1_QPLL_lock,
        s_axi_tx_tdata             => p1TxTDataUp,
        s_axi_tx_tvalid            => p1TxTValid,
        s_axi_tx_tready            => p1TxTReadyI,
        m_axi_rx_tdata             => p1RxTDataUp,
        m_axi_rx_tvalid            => p1RxTValidI,
        mmcm_not_locked            => dPort1_MCMM_NotLocked,
        drpaddr_in                 => lLane_DRP_AddrIn(1),
        drpdi_in                   => lLane_DRPDI_In(1),
        qpll_drpaddr_in            => (others => '0'),
        qpll_drpdi_in              => (others => '0'),
        drprdy_out                 => lLane_DRP_RdyOutSlv(1),
        drpen_in                   => lLane_DRP_EnInSlv(1),
        drpwe_in                   => lLane_DRP_WeInSlv(1),
        qpll_drprdy_out            => open,
        qpll_drpen_in              => '0',
        qpll_drpwe_in              => '0',
        drpdo_out                  => lLane_DRPDO_Out(1),
        qpll_drpdo_out             => open,
        init_clk                   => DerivedClk50,
        link_reset_out             => dPort1LinkResetOutI,
        gt_qpllclk_quad1_in        => Port1_QPLL_InClk,
        gt_qpllrefclk_quad1_in     => Port1_QPLL_RefInClk,
        gt_to_common_qpllreset_out => aPort1_QPLL_ResetOut,
        gt_qplllock_in             => aPort1_QPLL_LockIn,
        gt_qpllrefclklost_in       => dPort1_QPLL_RefClkLostIn,
        gt_rxcdrovrden_in          => '0',
        sys_reset_out              => p1SysResetOutI,
        reset_pb                   => dPort1CoreReset_pb
      );
    -- Reversing the Data Values
    p1TxTDataUp <= reverse(p1TxTData);
    p1RxTData   <= reverse(p1RxTDataUp);

  end block AuroraBlock;


  -------------------------- Unused Required Signals ---------------------------
  UnusedSignalsBlock : block
    -- Initialize unused signal so compiler won't optimize the signal away.
    signal dZero                    : std_logic := '1';
    signal Eth1GRefClk, CpriRefClk  : std_logic;

    -- The dont_touch attributes must be applied to the CELLs, and not the nets
    -- that are optimized away since they are not connected
    attribute dont_touch            : string;
    attribute dont_touch of Eth1GClkBuf   : label is "TRUE";
    attribute dont_touch of CpriRefClkBuf : label is "TRUE";
    --vhook_nowarn UnusedSignalsBlock/Eth1GRefClk
    --vhook_nowarn UnusedSignalsBlock/CpriRefClk

  begin

    --vhook   IBUFDS_GTE2   Eth1GClkBuf
    --vhook_a CLKCM_CFG     true
    --vhook_a CLKRCV_TRST   true
    --vhook_a CLKSWING_CFG  b"11"
    --vhook_a I             MGT_RefClk125MHz_p
    --vhook_a IB            MGT_RefClk125MHz_n
    --vhook_a O             Eth1GRefClk
    --vhook_a CEB           '1'
    --vhook_a ODIV2         open
    Eth1GClkBuf: IBUFDS_GTE2
      generic map (
        CLKCM_CFG    => true,   -- in  boolean := TRUE
        CLKRCV_TRST  => true,   -- in  boolean := TRUE
        CLKSWING_CFG => b"11")  -- in  bit_vector := "11"
      port map (
        O     => Eth1GRefClk,         -- out std_logic
        ODIV2 => open,                -- out std_logic
        CEB   => '1',                 -- in  std_logic
        I     => MGT_RefClk125MHz_p,  -- in  std_logic
        IB    => MGT_RefClk125MHz_n); -- in  std_logic

    -- Unused 1Gb MGT clock on the USRP RIO.

    -- Drive unused I2C lines to high impedance to allow board pulls to take over.
    Port0_SCL <= 'Z';
    Port0_SDA <= 'Z';
    Port1_SCL <= 'Z';
    Port1_SDA <= 'Z';
    --vhook_nowarn Port*S*


    -- To drive differential outputs, we need a flip-flop to drive the input of
    -- the OBUFDS. This flop is initialized to a '1' in the signal declaration above
    -- to keep the tools from optimizing it away.
    PackedFrag: process(DerivedClk50)
    begin
      if rising_edge(DerivedClk50) then
        dZero <= '0';
      end if;
    end process PackedFrag;

    -- Not supporting CPRI so don't need to drive the recovered clock to the PLL. To
    -- preserve the IOSTANDARD in the constraints file, we need a differential
    -- output buffer. Otherwise, the tools will complain (mainly just ISE, but possibly
    -- Vivado as well).
    CPRIObuf: OBUFDS
      port map (
        I            => dZero,
        O            => CPRI_RecoveredClkOut_p,
        OB           => CPRI_RecoveredClkOut_n
      );

    --vhook   IBUFDS_GTE2   CpriRefClkBuf
    --vhook_a CLKCM_CFG     true
    --vhook_a CLKRCV_TRST   true
    --vhook_a CLKSWING_CFG  b"11"
    --vhook_a I             MGT_CpriRefClk_p
    --vhook_a IB            MGT_CpriRefClk_n
    --vhook_a O             CpriRefClk
    --vhook_a CEB           '1'
    --vhook_a ODIV2         open
    CpriRefClkBuf: IBUFDS_GTE2
      generic map (
        CLKCM_CFG    => true,   -- in  boolean := TRUE
        CLKRCV_TRST  => true,   -- in  boolean := TRUE
        CLKSWING_CFG => b"11")  -- in  bit_vector := "11"
      port map (
        O     => CpriRefClk,        -- out std_logic
        ODIV2 => open,              -- out std_logic
        CEB   => '1',               -- in  std_logic
        I     => MGT_CpriRefClk_p,  -- in  std_logic
        IB    => MGT_CpriRefClk_n); -- in  std_logic

  end block UnusedSignalsBlock;

end rtl;
